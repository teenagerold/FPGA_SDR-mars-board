��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"a5���f���wR����.F�o!��5���?��Ԣ*5lkc�B|�yk�zzhT�1 �HAX��S�����jZ�w���EpM�\��q�sF'5����ɯ�@� ��@� �������ۄ��>���Յ��f�S8(/������a�M��ڗ�p>}�K9�� j!#����/��P��7c�p����꽈�ܼi�/�ǉH��S3��/d9Ex�~ ٢K�>����C�$�� ��=�D��Z���Ե��a�
��Sf1?U�c\��w��!�p��;nzY�~}��h�`҉Y�&�	�X/�>�����=��pu�~-y|TsLC0��i�1�I��x���SsA��;�񮗴5N	�oZS뛗�I{�r�s�JOOPZ����R��q�õ�N��WI���j9�����L[1:D���6�I�-~� oJ�L�Kz~:�# |b�咄t;���]��nM=
��C?������G=�R\V�"��S^8��ݱ�L���i��A���'��"�6�+��o��_/ ���:V7�5x�t�xg¥]���
w�Q.F��p���̠��M�V1D��MV�LS_Ҝ ���
��[��{�>M)n�
'���::GxeA��5
7Q�3Jpݗu$T��$�ދ(���w%��L�)=#�{����kJ6��	C�*+��B��p�X��c�{��b���ޭԐe���F��}���Z�:�	!�E!ϱ�#s����aIPL9\�$*���,�-J���y�3�k靯k�W��ȗY���Vq�9�s�~_<�2�'<��(0l@W��dά��ƿYZ�4�\z�ԺR3��+�V1_�O���[i��a{ᶸ�V���}V��5}�Rw������P2�"��똷����& T�)�_�}�	0keI���*}���\�z�B7 �)�m�4N3;�`�L�jQd&R��F��j�]x���n[�PӸ����y�ŹF_��J"ĭ�ѶF� ���\�;�ev����x�A��9���̜\�7��+5U"4Š�GQO�"@�T��n��3'n�|ב�]~c"O�ʛjL��p��H	�P�t8s�&$�-䷹DY<�*���r�ݎ孄w�%��dls���
c�������Ԍ����P��e�|�~���J:���5bEM�2K� ?�Hg����'Ȓ���އ�#����&�㭙1o�7�K���5��������P�E�y��J0ͧ-�{�l��C8��L�r��M�iڽ���:��	���v����7\����|	c`��5 V%�"y`.�kI�� ���B�?�?�,U�T3�4��&Č�I�d7����^�V4!3��y�>�D�383��������yC���E)����e�@-|���=�!_�5��`�ġ5N�����	p�@���niWKY��-7���%v.����3|�X��HN�Tk�I�`���	����GK�m�k�d�#MQ�n�cڎ��I7���H�,Ef�J4���<��&"��8��$rq�>���\���{X�^;S}�0��!z��t�{���|���r{�,�}�4�S,o@�
!E��%��v�@�]��ɸ��"��8ŕ�B���k�te�i�?��Ag�]Ճ�1"^֡�%�A���c�xg�E*<ܨڃ���\pԇ[\r�^��*u1������u��	�\�g���:zڧA���7(�B;:��_:���oh �Fk���_e�t3E"�<Q�V��	:/��^�4s߯ƞ!����j;`A'I�2E�V!E���(��ْ�ar���u%������Y3��u��ȿ1�OU����7!9�9?��E＀�
Dr�d���t<e����9G�����v�f�r'�����%-���U�'���lfZU���P��ϱ!��c�pf�9��Y���r�C���`
���l)�f_�hY�,%��������H��%56>��0��	��8�MSH~�1㸉����	�J�ck��7`1� �{�Pƶe��0�6��^M~N}5K����1rz��Mv�ԐiW(9.��2��f��ʒ
r7��F��T�6�j��x��hֶ۵m^u�ZT����N�\����X�~��@ ��q�����w���nbb��J%��\ꭊ��o⚰����!Nᑚ���O�����M':��V1	���BYsO~��J˨�1�J�sd!"�-O�<��5�:���{��Ž�z�zxy���ߚ����ҥCvtR�7�xf�g���
+V� \�6�R�Cy�_R��mf[>q�ʠ8
��ڌga���qd���>�K4q|9�Y�!ڕ��:�������@_�9�E�j?�G�{m�����(I��F��w6{��2�;1����oW.�"Zw��0���f�p[�Q��!v�Hz���f��W9B_̟��Y���M��i�>r�3���i��J �l>x#6	�K2l�~	�4�<�F� �N�V	��sp��CzAK�ת���r|�T��S�	& I��{q�k�+�ܶ ��D4'W�siRյ�07�X�8X����7�Md)�@��y`���u
���ٰ#�4z�A�j�|�/��0	�l|�J�B���Zy��Ek�,b��r@�����WG�v�<XO�!^�b����3ೡ�U�)2MQ�Kde�ߴ����Y��;���2ORR\���G9�~H?�fo�݇�L����s���?���=��O����$�i��k�#V��ɗL0 ;nd�7�$+b���=*N֢f+4V?����@��:�����t�z�>��zz2���`�{���3�������x;W�)nl�p��&>��{�"�aF�.�f��{�l��)k���{��)��w���3�i���6�#qh%��뿥���L��M�¥ŗ��l5�݄���WW��wﴌ0��)��u�9h�yy�L��[K�[/���r�k^b�n�u���u�ui�=���q_EXA:��!?��3�h��|߁I�'�����hq��7h�Q�a=��1`n�*��؋���A��c�8��탋�h��\{6�m~�g��[�ø��\^XPr�c����Zd^]�[�gv��"t�¸���WF����)�����_M&���46,X�K��t�����M� �ga��	���@8�?�qsBǨ��>��vҽZ���d]dU؍^%k��p�4S�6�o����+�Ho�SV����F���t�>V������5�C���{����n��:��B���,>�C�Z���b��obkB���P�Z/$�)��ڛ���jxϗkW1(�]R�y��Zy�<�[<3��r�	�a-����M��ў���xb���[�Z�M~�����-^�J���Z\0��i��ӡ]�lWe;#��4���R.�L��>�;�F��ˋD�L�k~7h_B|qAb�T	AÃ�%���uur$�wE�ʌ�C�t���6�4�l"b�ˡ	��jc8��@e��<�k]D�o��I�����ĺ�.oY���Ҋ�%��G�(�8�_��	W�\��JC3n���u aAm�;���0���@X.����S���*�S�T:fM��K��Z?5Y���L�._?����]�K*pl��D�B3(n���� �a-��x�aW�m���4��cL��U/E��3��kw�5��@���u6u6�K1���iN4��kLO!���o��s�]c�1����#.�Jrκz���4A ؜#jd	� ���4�j�q�U�5���ܲ;	Tgft`:�k��"��� yk���;�Z���}��Vz4�����3H)���B�J�Bݎpd��mȣ��p�����y�匿~��o�W쭛1S9 ����٨�$p�.��|�5� ��5<Gpԃ��W���I>�0M�/lY/br���4���^4:z��+������i��He��ʄg ��Ҍ�9x/�5;�Noт���������7���B���� <G�ѻ��z~������T���S������A�\d��޲��'�cy!����H�X5̅��E�~!~��]㿤�:h����d;��$����mbN{�tO��5Z�7ؤ5?Iq� �[:�YJ_;��*���:<�%��>pI��Z)��F�����ծ���aY���ņ:f�Y��V�ї�pb�;�9K��s#�d+<�H)bX�&��Q|��d�U��?��a���v����E۫_d֧�DM7S�օ��a�����J��s��o����X_{���ЧJ�Q�)�Ơ�b�`q��nb<gu`����*J��5�}��%���Y�������>8u����<���P�5��k��ĭ���b����z��Q�U��O�ma��X#�m(ÄR�~xfB:I�x����e_]}"(:�	�ۮ�8 ʑI�l��]TAY>s�򆼡���p�|�D)�m(�cu���p��'��|)������1���o3.]1\Dm�ϋ��)���1~���{��~��tt ��� ���9/��z�]��!񲂕��J�s汄#�Q.���cpՌ�C�8J
�F�V���l;}C�v�c�s��q
?���%�O����&�zy����?��O�A	A
�|���4�EmGº���1����ӧyW}�`;ul����h���2T�����/�1�SY��¶�u�z6�aL�s_�E0K��hHy��E���[g��@F|�MYmhl�� l^�l.�	E���LԴ<��Pe ����8��r�Þ)L	��3�6_�]0.^	f��C�PAe[)|��(-����]�U��j��yy)��GS�)�Ns��X��UP 1�!���PD��Q�2}O�{�x��3Lr f.����:͠�[�D@ڛhaP��:�؛h�D���-{��O���c��I�F����CE��Y�8�"ǂ����
�𠁕_ώ�P����!��@��#]�{O�<�HA�*��K��l�;�"��b|P6�a��. �dE�����6�����#�a؅Z����)]5BD���(��գG��A�Z$-��׭� r�9{�n#wA`�$�=?�5��1��e���G>�Y����+49N�$&��������B���F3�����B�q)�Y���to�A�1����:|��C��߲QO�^�v�.��넶g��`R#hAŷ��h_"�\�NE�9n�12�ӎ�Y��;�!ѧ"|�Y�iS�ȡ'vboo:7g���=���#�������w\Xk�k0]�|�fD�Z���h?��2̀�S�?%��R�)m���w�o��ᠫ�Ǌ�޶~���eV� 8�ZxN�~��I3ͽ�L��ܠ��4����E�����J��bƞ:��68���o.��1$�5��UB �i�&�R��(OKHki����JK�?�"���t�Ŀ�o��vA���[$��-��: �9�ÐK�η>=Dj��������'C�y
E��jF�[�-*y�]q��~��n�BMo��3B�(�O,����'���s�ɕ���� ���@D��ŠDa+��?A�"m�Ncp�l����蔙��m2�٣�xښ�%d�����ʺ�Ū8��K������<��N֤H#1���H�t��S����z����{��������	�ՒE ��A��?���k-J�t�U�-�z,�{~g����:��D%��i~�(��~�_���>�o�.ǧH��-��1�+Svt3\�K���1��Rsݏ����M�����4����YM�<�� H��a�����t�T�j���!�����d���u�@/g��M�H0T�l�09��0%fC2+�\�U&�jfב��5���J�»v�m�tͮ&9��	낳���~u�n�L��wsA��Ay�k_ �9��!�2���c�W������p~�n�l���R?����^�Ê3/R'K$s��b��6��*:�5mѷ����P%dW$�����׸�&i�L��n5[�]�Bq�!X/�'�Ν��l��.�ij�{����L ^���������E0��R��w;D���Z�gz��c����Q��P�g�={a.�{�yOC.;"�0e�G��u2��7�feW,]�"R9���x��S��;;K��l,��g/Q�a�iO�7�G �Lfʇ.�r�D�Îo{�vF]Y��'G���dA�u秘cI�'T��UQ�Z�݋�:�{���q�� b���D�M�N�rBE���^�E������n7������}���Η�9�U��.y�� �
'Yo��bk��e �%�]٠Z����81�������\�K����N�AXT�q�Mv�8��A����ч�?��.v�?٬wO�Iz��#D-�oAf���C���^e����6�q���h��X׼�ʝ�=�U��x�������&��\���a��6�[N�G��F�T�_��[ �u@�h9��J�v9��;���:=��*w�[��ŗs������vW;�Q"��Q���]/L�DS8v�r��6���[	z�zj"�@b�|�"εEgO�"���K'���5G~6�S���19[��"�	����:>����W����o��'ݔ�i� ���^h) ZxJ�^��n�y��vѿO6 ��v��W�.%ʼ��#wS���If�O{2��kѓdU�)f[��;�3�y��HB'}�>�a H�DBT���^� �8�"�5M��tq�5�<���9�畛��ϳ�������	��f��4W�ޒ$�����{7�9B+㹯�k�#��[�#w���uD~��|�H,�x���Yc�yBJ��;�����V��:���-qޥkW��2��q�)��s
��x�;�<ć8Thۙ�E�j)����$��&\*zi������i%,.�5�L�]���H��bk7y�?#,hz$/u��ø?��_�Y����k�iEd�U[��P�`?'(�3�7n�e�b�;{=c_�fJ��Ŭ��( q��W�L���l�2�Y�r�n�q"[?����r����!i$@���#��f�|�3%wI��C�a�jjD^�cW��j{S�4��$��M �Û�����/[����/��ܭ�K�Z�����Ks0�A�J �\��J�5�V�҆�z>x�N����@�Fx;�\I�#���$�y�z�ø(V��]���Kd,92��$[n��&`CL��N�5C�z�}�V�	���B��]4W�����[1;
\i�w��.3�L��X�~+�)A���}�h�m�-�(f�sʺ�I�ZJ�;w��^e W��W���5��F�&T�q��NQ0�F�Bҡ�EӸ�Kp�\�L;j�$�[4>hNF\>nR{Dl4�'�M��ʀc6�BP'������'�В"G�O��Ģ�N���5��(%����Қ��\WК��x>^����P=CKl?������ԭ�}(x�!I�}4�ĕ�%ɮ�Um�Y!���QJ���S��3��.z'Y�GOw'� ,#�29�&b� 2�W�;����nt�񺻟Ó@1���6���7[9B\f�`���G��R�[d���Ӱ�ŝ�n>0�'�8�Ԃ�}c}=lc��>C\h:���dd����X����O�f��ޜ�X����p�Lޮ_5�00p��8F�c���+�D�\���v�=��ٱ��Y��h��'��_A!�|;�g�W%̺=���gwګ��hY��g��#��f���,�	�����R�=��LD2�NϺ纆Z�8E_=���1�,K�w26�{���u9������eV�)!��ȕ[w�����[ZL�ʑ��<�^�p~lyDE�0Cs�wW�jEӧ?AԱ'�*�r���7{�H���W;�#�a:'w���r�q�w��2�g�OӢv~B�~���f��Q�¨O�����NY#����D�Wy���nޮ�t�Hr7�P�ZJ��־-s)��'bm-��A-�A;i�$�o��}I��2b�>n�1S�%����"ZY��P���g� ":�T��к
	oвH��x^�g�0º`<�5���ݲ��K�p�/��`$|�v�[*�ˈ��0�e#���V7������~Z�;V@8�-ؚS G$;�	�`װ|s�J�躖lt�H	h^R(&su3�
9J�ǆ2�a��D�~3���!+*I.���5�������&�o��s������>Z���*�x&d=*��I)I���j7��M%&|gY^�it�MʯkIH������o�N&�u�"�X�@��w'����2�~� :݀�Huu�-�!8\WN���=��f��oӓl��g�H��Qx�is�,f�b�!Q��Vt`D�A�O=�r���Wj���Hջ�B�ʗ�𛠳p#Wv��x�^������l�G�YGd�`M����_�=*��3�0�2��!���v"r_�4�1@}���u�ƶҞ��g_�8Y;������#����?{� �FB��E*�/z)��fNk��uPN�D�9�'F�WUr���%ɔ�^�V/3�L��\5,��a:���2��)�7k��Aӳ�3���=ت���.��	Ka�b!��6���[V�O�0�l><k[�r��Mۧ��g���log�(�]����^t<�\�wOS+Ut�%n�6�:�a�����Uh���T<���F���wu���flr�6���/>��!��l�U		�OZ)?_�#�Z��?OƠNF�J��K唾��GW��NA�+�B���U`����4GSHq�d,ϩW=�<�Nr�/���7��Va@"�k���������<���[9�TL��Y�W
*o�H�j�Y���$I�d;�z,WGOewK�B��Z xd2zf,/���w����	4	U4A�P΀9y�=�No�����>�k���gR!k	e�*���sx�Ey'*���+>;����~��1(�����zP�m��8�22����b�^k�p%p�?��t��K�C�t.��nql�*2
֣0'~Z&Ln"��,gp>�/c
+G��-��F�g�0��+o�ҫ���h�;��\V���b�������ZV�?��d��Z�0]�UU���-rP>��uv(P*�%:�$���-bI���n^�}�h�q,�	����~�[�}��]S����	��\癬��	�Q��
f�fG��ê�߮�}�܀�ie��F#-t�4�� r�k�tTon��2q#�]��pT\Ȥ�&��������r$�pr�&-�8��kHR������nN<��Ο��m.j!O�o��٭��e�Hwx���-����
���1:��u�\N㨤i��$|���Vk�(���)�;F�z�8N���lnV��$8[D򛏿W��4��Hy4�k�T�&�3?0� le�+����
�bbG���<Cb7���L�}�3�0.H:��i�����A�x�.{lָ� �I"y���?�@c��Ϣ�`Y�T5�?�P�ϯ�j��*�����h���QQV��B�PT�
�@)?.{����`�Y%��g�F���A4��gT���Y2���^ӫ�b5�¡t��i��/��a��7k��]��4&Sıvy1�~�"�0�d�`�9��Gl(�K���jy�옃�i�δ.�V9��,���*/�_?Y�&����`|���F*���K>��y�J���Z��H���X_VpE�8b��Hَ����0�ڮ�t8���co�~�_I[��E	5��!nُ�g4m�\��L_�������N���C#eߧW3u�=��P^ArE�(`��7�H�(����`�4v���P�䴽|���ڏ�38��eL0����Z�(1�!=)3MC���iZ�h��n�ɕ�qH�,�� ���:Е�B�w�s$P�ޟ]=���c�/,��0�O!�����wsn�}��m6�4�ś�{๐b��Sv\mÁ��˺��55�C��Z��fy���/���ҋ����l��-���<W�	^�fۇ
�W�U(L�3�7�"�M?sy���R���4����U��p3\��1xa��э�p�Ct,��~�[2�t ��y�dk�w#.�/���m"ۮ��qy�(�j��Üt���v�1�\�_B�ul{OU|/t��f���U_��c�СP\���pl�EMa��P�C�chq!��i4��7O�~l��{CQ���iC8����,�U�5�N/	�B%���^YNE�n�ݣ���uq�%��}-lX�k;�=0� �w�q���-�+�3ϒ^H
�X�h�t&�]�GI�ȡ��P��#��q������ZV�\o�T���Ln�X%��HCv3>ץ�̀[�R`|u�x�{X������t��v%8$�3���z �;a��ײa�4��&������SM��%AB*��G��dV`�.�;6U�Z)��#g6��pS�n��t;,���%��[ӃƦF�iF�{����!ڈ����Ś��h?��爔}��K�֮�K��cD���2��$6o���w��r}��=<�_��X$�(�q���)�<H��Sୢx����T*�FX�[]\g�����9��O5�@�39���U�)/���yU�b�Ĥ����۪�)`������5�<O[�e��*��W�@�y�Բ����J�����#�:7�V�}��t���)8P�I���#�El8�P���8���|;
��P�Ơ�C:�,�v��@�u��c`��+=�I�n�W���Fy�u���^z#B����D�7�^���;�i���z��B�YPg�<�����X��An�f���>� !9�������i�C�j.(�E���A�y]g"��6e�3)yc���x��4 �"�|rB� /h���R&�Ϻ��^�D�d>F6�Wan:H�����o�c��*��r�7r>��M��CV����(n6� v��+������]y�Eӌ��ӓg<^ľG���_Z��k���bg#�&�-��,M��>�&g�0���!HV��=E��NR.	�����g����ּ�+���1���F�#Z%�DL��`g+��[�x��\0(�WBk.��ׂy�M�|��W�9rCMY^ ˏ��6�&rY'|���7�-uҦ
��9c
�0���}]�u��\TO��m�m�㌐��&�]+-Zv���Υ|1c��|�`D�{��3���H���MP	���Z�+0�4vM��<���C�I�ZSx \H� ;�n+�DF���1�ݟ�.]�zȉ���g���)"8��ȹe���z��,�:W
]p �����Ԧ�A0�瓎�8�����s<~'�� ��tjN�}l�T)�`<�9eO~�p�Zl]��U 	�L�&�&�?ߧ]W��$I����vu�6��αwM���W��8�,���Y����:5��3��
{"�4'���
��«��V��!��,��r��]l��N@7)�ZB�:�����%d��j04�-3}���Ǘ��%5��*���P����2�΃��]e��cA1��Դ'
����C��5��Cqڃ�M�����vu/9SS�ԕ��r���J������gD��� <���ʹ���K�Ĉ|�����?�$%ἉC�o��)��4M�������m��8mՒC��2��(M��M^yA&�ٝ�)�=�
�� $��C��H��jc��@LUV��&eY�/�����ݦ�* ��2�'<V��.�W�,?��R���B�Z}G� ��Z.o�-� k��J�Y|U�M�F�� �d
��5�;~L��m�������c�� ���M��j���|��iCb�:F�\��|Dz����#9��z���8���`{5Q��A�7�y�v��OM�j�	����!��hg4��ʍ�'&@�o6�c�>�75�Ǧl?d����;b4�|c<��I����G�꾶��<�9�,ɲ6
�c>���Jý��z~�dX�_Ux��?�w>C�� &�F�?����1�H�H�G&�%���1O�k Hޔޔ��w����?±�R$e69EmW��,��6:�0�`�YRv���"��,�h
V7m�b�K���>���%���~^�N���aA|s!]g��]�$���%�IA���6��f�?���3ϸ	�����GQ�v��/�2�gR<~n��V�Bnve�A9��BdFS��i�@~��ضR��GL�ݠ�݃�c;���D>㤲V���M�j�aA[Έ�M�Џ��瞾�9�����@%$��|x}�ʡ9 �v���7���%���D(S����ߦg>6���bt1��s�؆6(���J�L����<�G0�����7�������r��ϡ.tz�1��H�E+&-����#f��H�D�%/Nr�Ӕ2ý/zY���>��K�i��\!�v�r���,����Nח1��p��U���I%��7rP��ˋ��z�i�w�п����d7R�-ۛ>�ȇ�/�#�p�+#+��r�X��$u��(8�K���SR��jiF-H|��tP�5�'��w�s�B��@B��N�eM�߲6˃c�Ս�q�q��|�� N��5�����Gj_��.e]V>J*5A�
E�QXq<^Nm�(���H>�U�DɶZ�k�1s�����L�_	�g���F�ΆٕX�q�}n�*,���亏�0�hL;-L�ӫ�)%�c�|[tiB�2��<{
�S��T�n'�웓#�R�V�$4 �	���I�'R֤9#K^����	���WI�F�f_?���-�/r<��|=�`��Z���T�ܪ�����%T5�k��������@�@p�j�2��͚cF��Y>�{����b_��oxX�NyzX[~��wf�W>��K�lHB�7ay��j跃ሱ��?.�*�`ի�7]��M�p�)@y�hs}�C�B����l�N�>l(F�9��U!w�vd�B>v� �G6�����l��8VRE�j�C¡
Jsf$��i�ܝ?S,k?澪&�,s*k��'��Z�&�&3��Ѵ��1b:�6e����#k�ULINVv(�{��|�¶�����5�H�:��9���YL�M3(̥� �qy����h�+x�%m� �����.F�V�j�8W낐��D�VBC^�?����/3��'i�k����K��@�`�M7�~���L���-�y �����ٶM���Q=ڷk�Ø���=�铣�d�����mhaK���#Vb���~S���[6INwnX$[�"��P�F�����:�@2	�,��1���ΰ]@R ���*\q��O���L�,	��2�JE!�V�hÊ��u�4 �xGVT�1�����iA��D�x=��4: ��Nz��'6m�^�Έ��YO�EN[Ss.�׌EC��t{vm�_T�y�����/�ن����������Q@�����[4}�F��rƳ�J8�5X`��(h��訔�����\GD[��j��LTQ�'�cL����fZ�4�%3)��~�2E ��i���:DI�{Dd��Hlb�UH�?�X?yO��Q��b�1�y
�^i)���-�ך�Ѓ}?t,1g��0��n�ܘK�1��1H>l���\�i�>˼qR'��2z����@��"���6'V)��de ��,����Ly0�L�)�`.�~����5�|���,@��3 m��t&i��c�#�B��?"V95˛Z%�d���)�c��$J�w�$�ݻ<į�Vrx�6

nz�.(�� E�b�<d��ĵ�����p��S�y���s¦�T�c�^K�W6�������n����"jn�$�t ������x�i!�`mآ'�s㯹���Oھ�xڰМ��Avp�m%��Q���B��H�����w�O���_��jH��D&#���� ����\��w?9���'mm�o�n	�u*Lz��ང��<f'�_�¦j�OzT���O�|!��n5)#�@�3�� k�mQ'K�Ľ�qx�m3x~9#ܶbo��&����4a��[q|D��2H�(��l�=�?n_qFG�G��Ƒ��/�z�}����R� ��'Sk�n�~g��/���uJ Vn���@����lM�걢�0�l�rԡ��(��f:P����s��]��j~ R�*�*���/��B	���e��u�7�JBAa��k����3Ǐ^���h;լ�m��kpm��j?:(�6�;�X��	��j:gs��Z�F'��/�li���7��;@s%�"CS��Z4�aGZ�nv�ư;r�4� ��XgP��*P�y�V<,�=��ZN�/�N>���,��3�l�*��"T���O�5��PO��|�"<H��D��X���%��|��a!�a�~v~w��
tׯ����3*���&���s��b���ᬞ��ܽ�86.��������q��*zb6�#�����B��6eMf���'���,��� k5? ��5p:�L�W8;�cN������U�ͺv�|Ap�K��O%e����S'c؏\-^��c
⑛��\�JD�ƨi"f?�l�X]:.�x~��f�͖��)�K�^o�������P��F�p��PcD5���0�Ga�k�(s�%ɛf�[�&� ��&�3�t�&ؒ��HE�'���rD�o�q��^d�I}y�G�Kr2*���R��Z�P1��G�[M7EAOBG���U���i>mk���8�4�c�ӛ����t}���SSg���Q��9_hs7�L!gf�����؄��n���F�|Q\a��lhA��k�ѭ]v�[q�7� B�o1�JyC
�%F*��ҔG�X�GTX�Q���K���kBSq$�@���ǭ*q�>+��Ҧ�����ԃ�@z|�i������6D�$@yR\�j���e�p/BS���	$�@�j�bz#�3K|��!b�M	H�F�E2%^�z�~�Vs��Bd|�YK����'�z3�i��:��L����b�H��U�PґP�O"� ��s^L��|c\�,�ٴߋV"��Q�9��ʇ���wF��5��k�YVRYDz5�.P5ؘ�O��zch+���/�~|U�$�o�f���}�)�HI�[3�"